`include "top_hvl.sv"
`include "interface.sv"
`include "driver.sv"
`include "monitor.sv"
`include "scoreboard.sv"
`include "agent.sv"
`include "coverage.sv"
//`include "assertions.sv"
`include "env.sv"



`include "test_basic.sv"
`include "test_int.sv"
`include "test_double.sv"
`include "test_dirigidos.sv"

`include "assertions.sv"